library IEEE;
use IEEE.std_logic_1164.all;  
use IEEE.numeric_std.all;     

package pRSP is

   type tDMEMarray is array(0 to 15) of std_logic_vector(7 downto 0);

end package;